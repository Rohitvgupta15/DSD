module or_21(
    input x,
    input y,
    output z
    );
    assign z= x|y;
endmodule
